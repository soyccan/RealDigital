module Compare(
);

endmodule
